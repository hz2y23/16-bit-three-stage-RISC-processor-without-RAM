// Wire widths
`define WORD_LEN 16
`define REG_FILE_ADDR_LEN 3
`define EXE_CMD_LEN 3
`define OP_CODE_LEN 4
`define INST_LEN 16
`define Gen_LEN 6

// Memory constants
`define DATA_MEM_SIZE 1024
`define INSTR_MEM_SIZE 1024
`define REG_FILE_SIZE 8
`define MEM_CELL_SIZE 8
