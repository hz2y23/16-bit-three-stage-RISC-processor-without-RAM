// To be used in side ALU
`define EXE_AND		3'b000
`define EXE_SUB 	3'b001
`define EXE_ADD 	3'b010
`define EXE_SLL 	3'b011
`define EXE_SRL 	3'b100
`define EXE_XOR		3'b101
`define EXE_OR		3'b110