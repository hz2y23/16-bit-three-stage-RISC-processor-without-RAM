// To be used inside controller.v
`define ADDI 	4'b0000
`define SUB 	4'b0001
`define ADD		4'b0010
`define BEQ 	4'b0011
`define BLT 	4'b0100
`define AND 	4'b0101
`define	SLL		4'b0110
`define SLLI 	4'b0111
`define	SRL		4'b1000
`define SRLI 	4'b1001
`define XOR		4'b1010
`define XORI	4'b1011
`define J 		4'b1100
`define OR 		4'b1101
`define ORI 	4'b1110
`define ANDI 	4'b1111